--4 bit binary adder--
--Declare library statements--
LIBRARY ieee;
USE ieee.std_logic_1164.all;

--Declare entity--
ENTITY lab2_1 IS
	PORT (A, B  : IN STD_LOGIC_VECTOR(3 downto 0);
			Cin : IN STD_LOGIC;
			 S  : OUT STD_LOGIC_VECTOR(3 downto 0);
			Cout: OUT STD_LOGIC
		  );
END lab2_1;

ARCHITECTURE structure OF lab2_1 IS

--declare signals--
	signal tmp1, tmp2, tmp3: STD_LOGIC;

	component fa is
	port (
		a,b,c : IN STD_LOGIC;
		co, s : OUT STD_LOGIC
	 );
	end component;
	
BEGIN
	fa0: fa
		port map(a=>A(0), b=>B(0), c=>Cin, co=>tmp1, s=>S(0));
	fa1: fa
		port map(a=>A(1), b=>B(1), c=>tmp1, co=>tmp2, s=>S(1));
	fa2: fa
		port map(a=>A(2), b=>B(2), c=>tmp2, co=>tmp3, s=>S(2));
	fa3: fa
		port map(a=>A(3), b=>B(3), c=>tmp3, co=>Cout, s=>S(3));
END structure;

--declare library again--
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fa IS
	PORT (a, b, c : in std_logic;
				co: out std_logic;
				s : out std_logic
		  );
END fa;

ARCHITECTURE fa_arch OF fa IS
BEGIN
	s <= a xor b xor c;
	co <= (a and b) or ((a xor b) and c);
END fa_arch;



		
	
	